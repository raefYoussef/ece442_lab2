library ieee;
use ieee.std_logic_1164.all;

package lab2_pkg is
-- subprogram declarations

-- type declarations
type char_array_t is array (integer range <>) of std_logic_vector(3 downto 0);

-- subtype declarations

-- constant declarations

-- signal declarations

-- variable declarations

-- file declarations

-- alias declarations

-- component declarations

-- attribute declarations

-- attribute specifications

-- disconnection specifications

-- use clauses

end package lab2_pkg;